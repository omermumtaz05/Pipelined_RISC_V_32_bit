module mem_to_reg_mux(



);



endmodule